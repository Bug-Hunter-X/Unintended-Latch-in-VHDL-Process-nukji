```vhdl
library ieee;
use ieee.std_logic_1164.all;

entity my_entity is
  port (
    clk : in std_logic;
    reset : in std_logic;
    data_in : in std_logic_vector(7 downto 0);
    data_out : out std_logic_vector(7 downto 0)
  );
end entity;

architecture behavioral of my_entity is
  signal internal_data : std_logic_vector(7 downto 0) := "00000000";
begin
  process (clk, reset)
  begin
    if reset = '1' then
      internal_data <= "00000000";
    elsif rising_edge(clk) then
      internal_data <= data_in;
    else
      internal_data <= internal_data; -- Added explicit assignment for the else case
    end if;
  end process;

  data_out <= internal_data;
end architecture;
```